
`ifndef   __type_defs__
  `define __type_defs__

typedef logic [31:0] array_32_bit[];

`endif

