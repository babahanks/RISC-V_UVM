`ifndef __risc_test_constants__
    `define __risc_test_constants__



`define  MEMORY_CODE_START_ADDR      0
`define  MEMORY_CODE_END_ADDR      100
`define  MEMORY_SIZE             65536

    // EDAPlayground has "Result reached the maximum of 5000 lines. Killing process."
    // So limiting to only 10 reg for now. otherwise 32

`define  REG_FILE_SIZE				7





`endif